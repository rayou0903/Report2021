----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:23:52 09/06/2019 
-- Design Name: 
-- Module Name:    top - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
Library UNISIM;
use UNISIM.vcomponents.all;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.ascii_pac.all;
use work.types.all;

entity top is
	port (
		CLK			: in		std_logic;
		WING_A		: out		std_logic_vector(16-1 downto 0);
		WING_B		: out		std_logic_vector(16-1 downto 0); --in -> out
		WING_C		: in		std_logic_vector(16-1 downto 0);
		RXD			: in		std_logic;
		TXD			: out 	std_logic := '1';
		DRAM_ADDR   : OUT		STD_LOGIC_VECTOR (12 downto 0);
		DRAM_BA     : OUT    STD_LOGIC_VECTOR (1 downto 0);
		DRAM_CAS_N  : OUT    STD_LOGIC;
		DRAM_CKE    : OUT    STD_LOGIC;
		DRAM_CLK    : OUT    STD_LOGIC;
		DRAM_CS_N   : OUT    STD_LOGIC;
		DRAM_DQ     : INOUT  STD_LOGIC_VECTOR(15 downto 0);
		DRAM_DQM    : OUT    STD_LOGIC_VECTOR(1 downto 0);
		DRAM_RAS_N  : OUT    STD_LOGIC;
		DRAM_WE_N   : OUT    STD_LOGIC;
		LED		: out		std_logic
	);
end top;

architecture Behavioral of top is
	-- ** component
	
	-- �N���b�N�W�F�l���[�^
	component clk_generator
		port (
			-- Clock in ports
			CLK_IN1           : in     std_logic;
			-- Clock out ports
			CLK_OUT2				 : out	 std_logic;
			CLK_OUT3				:	out	std_logic;
			CLK100          : out    std_logic
		);
	end component;
	
	-- RS232C�p�N���b�N�W�F�l���[�^
	component clk_gen_rs232c
		port (
			CLK_IN : in  STD_LOGIC;
			CLK9600 : out  STD_LOGIC;
			CLK115200 : out  STD_LOGIC);
	end component;
	
	-- �N���b�N�p10������
	component divider10
		port (
			CLK_IN  : in STD_LOGIC;
			CLK_OUT : out STD_LOGIC
		);
	end component;
	
	-- ��M���W���[��
	component receive
		port (
			RST			: in std_logic;
			CLK_RS232C	: in std_logic;
			RD_CLK		: in std_logic;
			RD_EN			: in std_logic;
			RXD			: in std_logic;
			FULL			: out std_logic;
			EMPTY			: out std_logic;
			ALMOST_EMPTY: out std_logic;
			VALID			: out std_logic;
			ACOUT			: out ascii
		);
	end component;
	
	-- ���M���W���[��
	component transfer
		port (
			RST			: in std_logic;
			CLK_RS232C	: in std_logic;
			WR_CLK		: in std_logic;
			WR_EN			: in std_logic;
			AC_TR			: in ascii;
			FULL			: out std_logic;
			EMPTY			: out std_logic;
			TXD			: out std_logic
		);
	end component;
	
	-- SDRAM�̐��䃂�W���[��
	component SDRAM_ctrl
		port (
			clk1	: in std_logic;
			rst	:	in		std_logic;
			--SDRAM�p�M��
			sdram_addr	:	out	std_logic_vector(11 downto 0);
			sdram_ba		:	out	std_logic_vector(1 downto 0);
			sdram_cs		:	out	std_logic;
			sdram_cke	:	out	std_logic;
			sdram_clk	:	out	std_logic;
			sdram_dq		:	inout	std_logic_vector(15 downto 0);
			sdram_dqm	:	out	std_logic_vector(1 downto 0);
			sdram_ras	:	out	std_logic;
			sdram_cas	:	out	std_logic;
			sdram_we		:	out	std_logic;
			
			data_in		:	in	std_logic_vector(63 downto 0);
			data_out		:	out	std_logic_vector(63 downto 0);
			req_read		:	in	std_logic;
			req_write	:	in	std_logic;
			address		:	in	std_logic_vector(19 downto 0);
			data_mask	:	in	std_logic_vector(1 downto 0);
			data_in_valid	: OUT		std_logic; -- �������݂�����������1�ɂȂ�M��
			data_out_valid : OUT		STD_LOGIC -- �ǂݏo��������������1�ɂȂ�M��
		);
	end component;
	
	-- sdram�ǂݏo�����W���[��
	component SDRAM_rd is
		port(
			clk : in std_logic;
			rst : in std_logic;
			
			rd_req : in std_logic;
			rd_fin : out std_logic;
			data_out : out std_logic_vector(63 downto 0);

			adr_in : in std_logic_vector(19 downto 0);
			
			sdr_req : out std_logic;
			sdr_adr : out std_logic_vector(19 downto 0);
			sdr_fin : in std_logic;
			sdr_data : in std_logic_vector(63 downto 0)
		);
	end component;
	
	-- sdram�������݃��W���[��
	component SDRAM_wr is
		port(
			clk : in std_logic;
			rst : in std_logic;
			
			wr_req : in std_logic;
			wr_fin	: out std_logic;
			
			data_in	: in std_logic_vector(64-1 downto 0);

			adr_in : in std_logic_vector(19 downto 0);
			
			sdr_req : out std_logic;
			sdr_adr : out std_logic_vector(19 downto 0);
			sdr_data : out std_logic_vector(63 downto 0)
		);
	end component;
	
	-- ��ԑJ�ڂ��s�����W���[��
	component state_machine
		generic (
			MAX_LEN					: positive := 64
		);
		port (
			CLK						: in std_logic;
			-- ��M�pFIFO�ւ̐M��
			REC_EMPTY				: in std_logic;
			REC_ALMOST_EMPTY		: in std_logic;
			REC_VALID				: in std_logic;
			REC_AC					: in ascii;
			REC_RD_EN				: out std_logic;
			
			-- �����񑗐M���W���[���p
			STR_FINISH				: in std_logic;
			STR_START				: out std_logic;
			STR						: out ascii_vector(0 to MAX_LEN-1);
			STR_LEN					: out integer;
			
			-- ���s���W���[���p
			EXE_FINISH				: in std_logic;
			EXE_START				: out std_logic;
			EXE_CMD					: out cmd_t;
			EXE_ADDR					: out std_logic_vector(20-1 downto 0);
			EXE_ADDR_FINISH		: out std_logic_vector(20-1 downto 0);
			EXE_DATA					: out std_logic_vector(64-1 downto 0);
			EXE_RESULT				: in ascii_vector(0 to MAX_LEN-1);
			EXE_RESULT_LEN			: in integer
		);
	end component;
	
	component signal_auth_ctrl
		port (
			CLK				: in std_logic;
			SEL				: in cmd_t; -- �I��p�M��
			-- ��ԑJ�ڃ��W���[������̐M��(0�ŃA�N�e�B�u)
			EXE_ADDR			: in std_logic_vector(20-1 downto 0);
			EXE_RD_REQ		: in std_logic;
			EXE_RD_FIN		: out std_logic;
			EXE_DATA			: out std_logic_vector(64-1 downto 0);
			-- ���胂�W���[������̐M��(1�ŃA�N�e�B�u)
			MSR_ADDR			: in std_logic_vector(20-1 downto 0);
			MSR_RD_REQ		: in std_logic;
			MSR_RD_FIN		: out std_logic;
			MSR_DATA			: out std_logic_vector(64-1 downto 0);
			-- SDRAM����󂯎��M��
			RD_FIN			: in std_logic;
			RD_DATA			: in std_logic_vector(64-1 downto 0);
			-- SDRAM�ǂݏo�����W���[���ɓn���A�h���X�A�f�[�^�A���N�G�X�g�M��
			RD_REQ			: out std_logic;
			RD_ADDR			: out std_logic_vector(20-1 downto 0)
		);
	end component;
	
	component command_execute
		port (
			CLK			: in std_logic;
			-- ���s�ɕK�v�ȐM��
			CMD_IN			: in cmd_t;
			ADDR_IN			: in std_logic_vector(20-1 downto 0);
			ADDR_FINISH_IN	: in std_logic_vector(20-1 downto 0);
			DATA_IN			: in std_logic_vector(64-1 downto 0);
			--** �e���W���[���Ƃ̒ʐM�ɕK�v�ȐM�� **
			-- �ǂݏo�����W���[��(sdram_rd)
			RD_ADDR			: out std_logic_vector(20-1 downto 0);
			RD_DATA			: in std_logic_vector(64-1 downto 0);
			RD_START			: out std_logic;
			RD_FINISH		: in std_logic;
			-- �������݃��W���[��(sdram_wr)
			WR_ADDR			: out std_logic_vector(20-1 downto 0);
			WR_DATA			: out std_logic_vector(64-1 downto 0);
			WR_START			: out std_logic;
			WR_FINISH		: in std_logic;
			-- ���胂�W���[��()
			MSR_ADDR_START	: out std_logic_vector(20-1 downto 0);
			MSR_ADDR_FINISH: out std_logic_vector(20-1 downto 0);
			MSR_DATA			: out std_logic_vector(64-1 downto 0);
			MSR_START		: out std_logic;
			MSR_FINISH		: in std_logic;
			-- ���Z�b�g
			RST_OP			: out std_logic;
			--** ���� **
			RESULT			: out ascii_vector(64-1 downto 0);
			RESULT_LEN		: out integer; -- ���s���ʂ̕�����
			EXE_START		: in std_logic;
			EXE_FINISH		: out std_logic
		);
	end component;
	
	-- ���胂�W���[��
	component just_measurement is
		port(
			clk : in std_logic;
			clk2 : in std_logic;
			rst : in std_logic;
			
			msr_start : in std_logic;
			msr_finish : out std_logic;
			str_adr : in std_logic_vector(19 downto 0);
			end_adr : in std_logic_vector(19 downto 0);
			
			sdr_req : out std_logic;
			sdr_fin : in std_logic;
			ctrl_data : in std_logic_vector(63 downto 0);
			cite_addr : out std_logic_vector(19 downto 0);
			
			test_dout : out std_logic_vector(63 downto 0);
			test_bit : out std_logic; --�e�X�g�p1bit�M��
			
			measure_output	: out std_logic_vector(15 downto 0);
			rf_pulse : out std_logic_vector(2 downto 0);
--			data1 : out std_logic; --DDS�E�p�E�M�E��E�
--			fqud1 : out std_logic;
--			reset1 : out std_logic;
--			w_clk1 : out std_logic;
--			data2 : out std_logic; --DDS�E�p�E�M�E��E�
--			fqud2 : out std_logic;
--			reset2 : out std_logic;
--			w_clk2 : out std_logic;
			adc_sig : out std_logic_vector(2 downto 0);
			IO_RESET1 : out std_logic;  --DDS3
			RESET1  : out std_logic;
			SCLK1   : out std_logic;
			SDIO1   : out std_logic;
			CS1     : out std_logic;
			IO_UPDATE1  : out std_logic;
			PSEL1   : out std_logic_vector(2 downto 0);
			IO_RESET2 : out std_logic;  --DDS4
			RESET2  : out std_logic;
			SCLK2   : out std_logic;
			SDIO2   : out std_logic;
			CS2     : out std_logic;
			IO_UPDATE2  : out std_logic;
			PSEL2   : out std_logic_vector(2 downto 0)
		);
	end component;
	
	-- �����񑗐M���W���[��
	component string_send
		generic (
			MAX_LEN : integer := 64
		);
		port (
			CLK		: in std_logic;
			STR		: in ascii_vector(0 to MAX_LEN-1);
			LEN		: in integer;
			START		: in std_logic;
			AC_OUT	: out ascii;
			WR_REQ	: out std_logic;
			FINISH	: out std_logic
		);
	end component;
	
	component vector_mux
		generic (
			SIGNAL_NUM	: positive	:= 64
		);
		port (
			SEL					: in std_logic;
			LOW_ACTIVE_SIG		: in std_logic_vector(SIGNAL_NUM-1 downto 0);
			HIGH_ACTIVE_SIG	: in std_logic_vector(SIGNAL_NUM-1 downto 0);
			OUT_SIG				: out std_logic_vector(SIGNAL_NUM-1 downto 0)
		);
	end component;

	-- ** signal
	
	-- clk
	signal clk100		: std_logic;
	signal clk100_nb	: std_logic;
	signal clk30		: std_logic;
	signal clk_rs232c	: std_logic; -- RS232C�ʐM�ɍ��킹���N���b�N�M��
	signal clk10      : std_logic;
	
	-- led
	signal led_inner	: std_logic := '0';
	
	-- buf
	signal outer_clk_buf		: std_logic; -- IBUFG, RS232C�Ή��̎��g������͂��邽�߂̃o�b�t�@
	signal rxd_buf		: std_logic; -- IBUFG
	signal txd_buf		: std_logic := '1'; -- OBUF
	
	-- receive
	signal rc_fifo_rst				: std_logic;
	signal rc_fifo_empty				: std_logic;
	signal rc_fifo_almost_empty	: std_logic;
	signal rc_fifo_full				: std_logic;
	signal rc_fifo_valid				: std_logic;
	signal rc_rd_en					: std_logic;
	signal rc_ac						: ascii; -- ��M�p�M��
	
	-- transfer
	signal tr_fifo_rst	: std_logic;
	signal tr_fifo_empty	: std_logic;
	signal tr_fifo_full	: std_logic;
	signal tr_wr_en		: std_logic;
	signal tr_ac			: ascii; -- ���M�p�M��
	
	-- crlf���ϑ����ꂽ��1�ƂȂ�M��
	signal crlf_observed	: std_logic;
	
	-- sdram ctrl
	-- common
	signal sdram_addr		: std_logic_vector(20-1 downto 0);
	signal rw_addr_sel	: std_logic;
	-- read
	signal sdram_r_data	: std_logic_vector(64-1 downto 0);
	signal sdram_r_addr	: std_logic_vector(20-1 downto 0);
	signal sdram_r_req	: std_logic;
	signal sdram_r_fin	: std_logic;
	-- write
	signal sdram_w_data	: std_logic_vector(64-1 downto 0);
	signal sdram_w_addr	: std_logic_vector(20-1 downto 0);
	signal sdram_w_req	: std_logic;
	signal sdram_w_fin	: std_logic;
	
	-- sdram read
	signal rd_fin	: std_logic;
	signal rd_data	: std_logic_vector(64-1 downto 0);
	signal rd_req	: std_logic;
	signal rd_addr	: std_logic_vector(20-1 downto 0);
	
	
	-- state machine
	signal rst_op			: std_logic := '0';
	
	-- execute
	signal exe_cmd					: cmd_t;
	signal exe_start				: std_logic;
	signal exe_finish				: std_logic := '1';
	signal exe_addr_in			: std_logic_vector(20-1 downto 0);
	signal exe_addr_finish_in	: std_logic_vector(20-1 downto 0);
	signal exe_data_in			: std_logic_vector(64-1 downto 0);
	signal exe_rd_addr			: std_logic_vector(20-1 downto 0);
	signal exe_rd_data			: std_logic_vector(64-1 downto 0);
	signal exe_rd_start			: std_logic;
	signal exe_rd_finish			: std_logic;
	-- result
	signal exe_result			: ascii_vector(0 to 64-1);
	signal exe_result_len	: integer;
	-- sdram write
	signal exe_wr_fin		: std_logic;
	signal exe_wr_data	: std_logic_vector(64-1 downto 0);
	signal exe_wr_req		: std_logic;
	signal exe_wr_addr	: std_logic_vector(20-1 downto 0);
	
	-- measure part
	signal msr_addr_start	: std_logic_vector(20-1 downto 0);
	signal msr_addr_finish	: std_logic_vector(20-1 downto 0);
	signal msr_data			: std_logic_vector(64-1 downto 0);
	signal msr_start			: std_logic;
	signal msr_finish			: std_logic;
	signal msr_rd_req	 		: std_logic;
	signal msr_rd_fin			: std_logic;
	signal msr_rd_data		: std_logic_vector(64-1 downto 0);
	signal msr_rd_addr		: std_logic_vector(20-1 downto 0);
	signal msr_rf_pulse		: std_logic_vector(2 downto 0);
	signal msr_adc_sig		: std_logic_vector(2 downto 0);
	signal msr_test_bit		: std_logic;
	signal msr_test_dout		: std_logic_vector(63 downto 0);
	signal msr_wing_a			: std_logic_vector(15 downto 0);
	signal dds_data			: std_logic;
	signal dds_fqud			: std_logic;
   signal dds_wclk1			: std_logic;
	signal dds_reset			: std_logic;
	
	-- string send
	signal str			: ascii_vector(0 to 64-1);
	signal str_len		: integer;
	signal str_start	: std_logic;
	signal str_finish	: std_logic;
	signal str_wr_req	: std_logic;
	
	--dds1 signal
	signal cs_inner        : std_logic;
	signal ps_inner        : std_logic_vector(2 downto 0);
	signal io_update_inner : std_logic;
	signal sdio_inner      : std_logic;
	signal sclk_inner      : std_logic;
	
begin
	-- ** port map
	
   -- IBUF: Single-ended Input Buffer
   --       Spartan-6
   -- Xilinx HDL Language Template, version 14.7
   
   IBUF_rs232c_clk : IBUFG
   generic map (
      IBUF_LOW_PWR => TRUE, -- Low power (TRUE) vs. performance (FALSE) setting for referenced I/O standards
      IOSTANDARD => "LVTTL")
   port map (
      O => outer_clk_buf,-- Buffer output
      I => WING_C(0)      -- Buffer input (connect directly to top-level port)
   );
	
	
	IBUF_rxd : IBUF
   generic map (
      IBUF_LOW_PWR => TRUE, -- Low power (TRUE) vs. performance (FALSE) setting for referenced I/O standards
      IOSTANDARD => "LVTTL")
   port map (
      O => rxd_buf,     -- Buffer output
      I => RXD      -- Buffer input (connect directly to top-level port)
   );
  
   -- End of IBUF_inst instantiation
	
	-- OBUF: Single-ended Output Buffer
   --       Spartan-6
   -- Xilinx HDL Language Template, version 14.7
   
   OBUF_txd : OBUF
   generic map (
      DRIVE => 8,
      IOSTANDARD => "LVTTL",
      SLEW => "SLOW")
   port map (
      O => TXD,     -- Buffer output (connect directly to top-level port)
      I => txd_buf      -- Buffer input 
   );
  
   -- End of OBUF_inst instantiation
	
	-- BUFG: Global Clock Buffer
   --       Spartan-6
   -- Xilinx HDL Language Template, version 14.7

--   BUFG_inst : BUFG
--   port map (
--      O => WING_A(13), -- 1-bit output: Clock buffer output
--      I => clk30  -- 1-bit input: Clock buffer input
--   );
	
	-- C0����̓��͂�RS232C�p�̃N���b�N�Ƃ��Ďg��
	rs232c_clk_gen : clk_gen_rs232c
		port map (
			CLK_IN => outer_clk_buf,
			CLK9600 => clk_rs232c,
			CLK115200 => open
	);
	
	-- �����N���b�N100MHz�𐶐�
	clk_gen : clk_generator
		port map (
			CLK_IN1 => CLK,
			CLK_OUT2 => clk30,      --10MHz
			CLK_OUT3 => clk100_nb,  --50MHz
			CLK100 => clk100        --100MHz
	);
	
	-- �N���b�N�p10������
	div10 : divider10
		port map (
			CLK_IN  => clk30,  --10MHz
			CLK_OUT => clk10  --1MHz
		);
	
	-- receive
	rc : receive
		port map(
			RST => rc_fifo_rst,
			CLK_RS232C => clk_rs232c,
			RD_CLK => clk100,
			RD_EN => rc_rd_en,
			ACOUT => rc_ac,
			FULL => rc_fifo_full,
			EMPTY => rc_fifo_empty,
			ALMOST_EMPTY => rc_fifo_almost_empty,
			VALID => rc_fifo_valid,
			RXD => rxd_buf
	);
	
	-- transfer
	tr : transfer
		port map (
			RST => tr_fifo_rst,
			CLK_RS232C => clk_rs232c,
			WR_CLK => clk100,
			AC_TR => tr_ac,
			WR_EN => tr_wr_en,
			FULL => tr_fifo_full,
			EMPTY => tr_fifo_empty,
			TXD => txd_buf
	);
	
	-- SDRAM����
	sdram : SDRAM_ctrl
		port map (
			clk1 => clk100,
			rst => rst_op,
			sdram_addr => DRAM_ADDR(11 downto 0),
			sdram_ba => DRAM_BA,
			sdram_cs => DRAM_CS_N,
			sdram_cke => DRAM_CKE,
			sdram_clk => DRAM_CLK,
			sdram_dq => DRAM_DQ,
			sdram_dqm => DRAM_DQM,
			sdram_ras => DRAM_RAS_N,
			sdram_cas => DRAM_CAS_N,
			sdram_we => DRAM_WE_N,
			data_in => sdram_w_data,
			data_out => sdram_r_data,
			req_read => sdram_r_req,
			req_write => sdram_w_req,
			address => sdram_addr,
			data_mask => "11",
			data_in_valid => sdram_w_fin,
			data_out_valid => sdram_r_fin
	);
	
	-- sdram read
	read_sec : sdram_rd
		port map(
			clk => clk100,
			rst => rst_op,
			rd_req => rd_req,
			rd_fin => rd_fin,
			data_out => rd_data,
			adr_in => rd_addr,
			sdr_req => sdram_r_req,
			sdr_adr => sdram_r_addr,
			sdr_fin => sdram_r_fin,
			sdr_data => sdram_r_data
	);
	
	-- sdram write
	write_sec : sdram_wr
		port map(
			clk => clk100,
			rst => rst_op,
			wr_req => exe_wr_req,
			wr_fin => exe_wr_fin,
			data_in => exe_wr_data,
			adr_in => exe_wr_addr,
			sdr_req => sdram_w_req,
			sdr_adr => sdram_w_addr,
			sdr_data => sdram_w_data
	);
	
	-- state machine
	st_machine : state_machine
		port map (
			CLK => clk100,
			REC_EMPTY => rc_fifo_empty,
			REC_ALMOST_EMPTY => rc_fifo_almost_empty,
			REC_VALID => rc_fifo_valid,
			REC_AC => rc_ac,
			REC_RD_EN => rc_rd_en,
			STR_FINISH => str_finish,
			STR_START => str_start,
			STR => str,
			STR_LEN => str_len,
			EXE_FINISH => exe_finish,
			EXE_START => exe_start,
			EXE_CMD => exe_cmd,
			EXE_ADDR => exe_addr_in,
			EXE_ADDR_FINISH => exe_addr_finish_in,
			EXE_DATA => exe_data_in,
			EXE_RESULT => exe_result,
			EXE_RESULT_LEN => exe_result_len
	);
	
	-- �M���̌������Ǘ����郂�W���[��
	sig_auth_ctrl : signal_auth_ctrl
		port map (
			CLK => clk100,
			SEL => exe_cmd,
			-- ��ԑJ�ڃ��W���[������̐M��(0�ŃA�N�e�B�u)
			EXE_ADDR => exe_rd_addr,
			EXE_RD_REQ => exe_rd_start,
			EXE_RD_FIN => exe_rd_finish,
			EXE_DATA => exe_rd_data,
			-- ���胂�W���[������̐M��(1�ŃA�N�e�B�u)
			MSR_ADDR => msr_rd_addr,
			MSR_RD_REQ => msr_rd_req,
			MSR_RD_FIN => msr_rd_fin,
			MSR_DATA => msr_rd_data,
			-- SDRAM����󂯎��M��
			RD_FIN => rd_fin,
			RD_DATA => rd_data,
			-- SDRAM�ǂݏo�����W���[���ɓn���A�h���X�A���N�G�X�g�M��
			RD_REQ => rd_req,
			RD_ADDR => rd_addr
	);
	
	-- command execute
	cmd_exe : command_execute
		port map (
			CLK => clk100,
			-- ���s�ɕK�v�ȐM��
			CMD_IN => exe_cmd,
			ADDR_IN => exe_addr_in,
			ADDR_FINISH_IN => exe_addr_finish_in,
			DATA_IN => exe_data_in,
			--** �e���W���[���Ƃ̒ʐM�ɕK�v�ȐM�� **
			-- �ǂݏo�����W���[��(sdram_rd)
			RD_ADDR => exe_rd_addr,
			RD_DATA => exe_rd_data,
			RD_START => exe_rd_start,
			RD_FINISH => exe_rd_finish,
			-- �������݃��W���[��(sdram_wr)
			WR_ADDR => exe_wr_addr,
			WR_DATA => exe_wr_data,
			WR_START => exe_wr_req,
			WR_FINISH => exe_wr_fin,
			-- ���胂�W���[��()
			MSR_ADDR_START => msr_addr_start,
			MSR_ADDR_FINISH => msr_addr_finish,
			MSR_DATA => msr_data,
			MSR_START => msr_start,
			MSR_FINISH => msr_finish,
			-- ���Z�b�g
			RST_OP => rst_op,
			--** ���� **
			RESULT => exe_result,
			RESULT_LEN => exe_result_len,
			EXE_START => exe_start,
			EXE_FINISH => exe_finish
	);
	
	-- measurement module
	measure : just_measurement 
		port map(
			clk => clk100,      --100MHz
			clk2 => clk10,      --1MHz
			rst => rst_op,
			msr_start => msr_start,
			msr_finish => msr_finish,
			str_adr => msr_addr_start,
			end_adr => msr_addr_finish,
			sdr_req => msr_rd_req,
			sdr_fin => msr_rd_fin,
			ctrl_data => msr_rd_data,
			cite_addr => msr_rd_addr,
			test_dout => msr_test_dout,
			test_bit => msr_test_bit,
			measure_output => msr_wing_a,
			rf_pulse => msr_rf_pulse,
--			data1 => WING_A(3),
--			fqud1=> WING_A(6),
--			reset1 => WING_A(0),
--			w_clk1 => WING_A(2),
--			data2 => WING_A(7),
--			fqud2 => WING_A(5),
--			reset2 => WING_A(4),
--			w_clk2 => WING_A(1),
			adc_sig  => msr_adc_sig,
			IO_RESET1 => WING_A(0),  --DDS3
			RESET1   => WING_A(1),
			CS1        => cs_inner,
			PSEL1(0)   => ps_inner(0),
			PSEL1(1)   => ps_inner(1),
			PSEL1(2)   => ps_inner(2),
			IO_UPDATE1 => io_update_inner,
			SDIO1      => sdio_inner,
			SCLK1      => sclk_inner,
			IO_RESET2  => WING_B(15),  --DDS4
			RESET2     => WING_B(14),
			CS2        => WING_B(13),
			PSEL2(0)   => WING_B(12),
			PSEL2(1)   => WING_B(11),
			PSEL2(2)   => WING_B(10),
			IO_UPDATE2 => WING_B(9),
			SDIO2      => WING_B(8),
			SCLK2      => WING_B(7)
	);
	
	-- string sender
	str_send : string_send
		port map (
			CLK => clk100,
			STR => str,
			LEN => str_len,
			START => str_start,
			AC_OUT => tr_ac,
			WR_REQ => tr_wr_en,
			FINISH => str_finish
	);
	
	-- write or read selector
	mux_rw_addr	: vector_mux
		generic map(
			SIGNAL_NUM => 20
		)
		port map (
			SEL => rw_addr_sel,
			LOW_ACTIVE_SIG => sdram_r_addr,
			HIGH_ACTIVE_SIG => sdram_w_addr,
			OUT_SIG => sdram_addr
	);
	
	-- ** signal assignment
	LED <= msr_wing_a(15);
	WING_A(2)           <= cs_inner;
	WING_A(5 downto 3)  <= ps_inner;
	WING_A(6)           <= io_update_inner;
	WING_A(7)           <= sdio_inner;
	WING_A(8)           <= sclk_inner;
	WING_A(14 downto 9) <= msr_wing_a(5 downto 0);
	WING_A(15)          <= clk30;
	
	WING_B(6)          <= cs_inner;
	WING_B(5 downto 3) <= ps_inner;
	WING_B(2)          <= io_update_inner;
	WING_B(1)          <= sdio_inner;
	WING_B(0)          <= sclk_inner;
	--WING_A(13) <= clk30;  --�ꎞ��~
	--WING_A(15 downto 14) <= msr_wing_a(6 downto 5);  --�ꎞ��~
--	WING_A(13) <= dds_fqud;
--	WING_A(12) <= dds_reset;
--	WING_A(14) <= dds_wclk1;
--	WING_A <= msr_test_dout(15 downto 0);
--	WING_A(15 downto 0) <= msr_wing_a(15 downto 0);
	DRAM_ADDR(12) <= '0';

	-- ** process
	-- test
--	process(clk100)
--	begin
--		if rising_edge(clk100) then
--			if msr_adc_sig = '1' then
--				led_inner <= not led_inner;
--			end if;
--		end if;
--	end process;
	
	
	-- read and write select signal
	process(exe_cmd)
	begin
		if exe_cmd = sdr1 then
			rw_addr_sel <= '0';
		elsif exe_cmd = sdw1 then
			rw_addr_sel <= '1';
		elsif exe_cmd = reqr then
			rw_addr_sel <= '0';
		else
			rw_addr_sel <= '0';
		end if;
	end process;
	
end Behavioral;